------------------------------------------------------------------------------/
--$Date: 2016/09/12 08:41:01 $
--$RCSfile: rx_sync.vhd,v $
--$Revision: 1.1 $
------------------------------------------------------------------------------/
--   ____  ____ 
--  /   /\/   / 
-- /___/  \  /    Vendor: Xilinx 
-- \   \   \/     Version : 1.5
--  \   \         Application : RocketIO GTX Wizard 
--  /   /         Filename : rx_sync.vhd
-- /___/   /\     Timestamp : 
-- \   \  /  \ 
--  \___\/\___\ 
--
--
-- Module RX_SYNC
-- Generated by Xilinx RocketIO GTX Wizard

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

entity RX_SYNC is
port
(
    RXENPMAPHASEALIGN   :   out   std_logic;              
    RXPMASETPHASE       :   out   std_logic;              
    SYNC_DONE           :   out   std_logic;              
    USER_CLK            :   in    std_logic;               
    RESET               :   in    std_logic           

);

    attribute X_CORE_INFO : string;
    attribute X_CORE_INFO of RX_SYNC : entity is "gtxwizard_v1_5, Coregen v10.1_ip3";

end RX_SYNC;

architecture RTL of RX_SYNC is
--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;

--*******************************Register Declarations************************

    signal   begin_r               :   std_logic;
    signal   phase_align_r         :   std_logic;
    signal   ready_r               :   std_logic;
    signal   sync_counter_r        :   unsigned(5 downto 0);
    signal   sync_done_count_r     :   unsigned(2 downto 0); --counter for iterations, for synthesis (5 downto 0), for simulation (2 downto 0)
    signal   wait_after_sync_r     :   std_logic;
    signal   wait_before_sync_r    :   unsigned(10 downto 0);
    signal   wait_stable_r         :   std_logic;
    
--*******************************Wire Declarations****************************
    
    signal   count_32_complete_r   :   std_logic;
    signal   count_1024_complete_r  :   std_logic;
    signal   next_phase_align_c    :   std_logic;
    signal   next_ready_c          :   std_logic;
    signal   next_wait_after_sync_c:   std_logic;
    signal   next_wait_stable_c    :   std_logic;
    signal   sync_32_times_done_r  :   std_logic;

begin
--*******************************Main Body of Code****************************

    --________________________________ State machine __________________________    
    -- This state machine manages the phase alingment procedure of the GTX on the
    -- receive side.The module is held in reset till the usrclk source is stable.
    -- In the case of buffer bypass where the rxrecclk is used to clock the usrclks,
    -- the usrclk stable indication is given the dcm_locked signal if a DCM is used.
    -- Once the dcm_lock is asserted, state machine goes into the wait_stable_r
    -- for 1024 cycles to allow some time to ensure the pll is stable. After this, 
    -- it goes into the phase_align_r state where the phase alignment procedure is 
    -- executed. This involves asserting the RXPMASETPHASE for 32 clock cycles.After
    -- the port is deasserted, the state machine goes into a wait state for 1024 cycles.
    -- This procedure is repeated 32 times.
    
    -- State registers
    process( USER_CLK )
    begin
        if(USER_CLK'event and USER_CLK = '1') then
            if(RESET='1') then
                begin_r           <=  '1' after DLY;
                wait_stable_r     <=  '0' after DLY;
                phase_align_r     <=  '0' after DLY;
                wait_after_sync_r <=  '0' after DLY;
                ready_r           <=  '0' after DLY;
            else
                begin_r           <=  '0' after DLY;
                wait_stable_r      <=  next_wait_stable_c after DLY;
                phase_align_r      <=  next_phase_align_c after DLY;
                wait_after_sync_r  <=  next_wait_after_sync_c after DLY;
                ready_r            <=  next_ready_c after DLY;
            end if;
        end if;
    end process;

    -- Next state logic
    next_wait_stable_c      <=   begin_r or
                                 (wait_stable_r and  not count_1024_complete_r);
                                        
    next_phase_align_c      <=   (wait_stable_r and count_1024_complete_r) or
                                 (phase_align_r and not count_32_complete_r) or
                                 (wait_after_sync_r and count_1024_complete_r and not sync_32_times_done_r);
                                        

    next_wait_after_sync_c  <=   (phase_align_r and count_32_complete_r) or
                                 (wait_after_sync_r and not count_1024_complete_r);

    next_ready_c            <=   (wait_after_sync_r and count_1024_complete_r and sync_32_times_done_r) or
                                 ready_r;


    --_________ Counter for to wait for pll to be stable before sync __________
    process( USER_CLK )
    begin
        if(USER_CLK'event and USER_CLK = '1') then
            if ((wait_stable_r='0') and (wait_after_sync_r='0')) then
                wait_before_sync_r <= (others=>'0') after DLY;
            else
                wait_before_sync_r <= wait_before_sync_r + 1 after DLY;
            end if;
        end if;
    end process;

    count_1024_complete_r <= wait_before_sync_r(10);

    --_______________ Counter for holding SYNC for SYNC_CYCLES ________________
    process( USER_CLK )
    begin
        if(USER_CLK'event and USER_CLK = '1') then
            if (phase_align_r='0') then
                sync_counter_r <= (others=>'0') after DLY;
            else
                sync_counter_r <= sync_counter_r + 1 after DLY;
            end if;
        end if;
    end process;

    count_32_complete_r <= sync_counter_r(5);

    --__________ Counter for counting number of times sync is done ____________
    process( USER_CLK )
    begin
        if(USER_CLK'event and USER_CLK = '1') then
            if (RESET='1') then
                sync_done_count_r <= (others=>'0') after DLY;
            elsif(count_1024_complete_r ='1') then
                sync_done_count_r <= sync_done_count_r + 1 after DLY;
            end if;
        end if;
    end process;

    sync_32_times_done_r <= sync_done_count_r(sync_done_count_r'high);

    --_______________ Assign the phase align ports into the GTX _______________

    RXENPMAPHASEALIGN    <=  not begin_r;
    RXPMASETPHASE        <=  phase_align_r;

    --_______________________ Assign the sync_done port _______________________
    
    SYNC_DONE <= ready_r;
    
    
end RTL;
